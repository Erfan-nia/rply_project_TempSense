cicsimgen tran

*Nothing here

.lib  "/home/erfana/eda/pdks/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice" fs

.lib "../../../tech/ngspice/temperature.spi" Tl

.lib "../../../tech/ngspice/supply.spi" Vl


*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../work/xsch/RPLY_PROJECT.spice

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

*.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
*VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VDD VDD VSS dc 2
.dc	temp    -40     125     5
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD VSS VREF VAMP V V1 VREF V-V1 RPLY_PROJECT

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

.save v(VDD) v(VSS) v(vref) v(V-V1) v(VAMP) v(V) v(V1) v(VREF) 

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100p 2n 0

*tran 10p 10n 1p
dc TEMP -40 125 5
write
quit

.endc

.end

